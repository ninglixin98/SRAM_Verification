`ifndef NLX_SRAM_ELEMENT_SEQUENCES_SVH
`define NLX_SRAM_ELEMENT_SEQUENCES_SVH

`include "nlx_sram_base_element_sequence.sv"
`include "nlx_sram_single_read_seq.sv"
`include "nlx_sram_single_write_seq.sv"

`endif//nlx_sram_ELEMENT_SEQUENCES_SVH
