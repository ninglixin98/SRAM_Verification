`ifndef NLX_SRAM_SEQ_LIB_SVH
`define NLX_SRAM_SEQ_LIB_SVH

`include "nlx_sram_element_sequences.svh"
`include "nlx_sram_base_virtual_sequence.sv"
`include "nlx_sram_smoke_virt_seq.sv"
`include "nlx_sram_diff_byteline_virt_seq.sv"
`include "nlx_sram_chipsel_virt_seq.sv"
`include "nlx_sram_rstn_virt_seq.sv"
`include "nlx_sram_illegal_addr_virt_seq.sv"

`endif//nlx_sram_SEQ_LIB_SVH

