`ifndef SRAM_SEQUENCE_LIB_SVH
`define SRAM_SEQUENCE_LIB_SVH

`include "sram_base_sequence.sv"
`include "sram_master_single_trans.sv"

`endif//sram_SEQUENCE_LIB_SVH

