`ifndef NLX_SRAM_TESTS_SVH
`define NLX_SRAM_TESTS_SVH

`include "nlx_sram_base_test.sv"
`include "nlx_sram_smoke_test.sv"
`include "nlx_sram_diff_byteline_test.sv"
`include "nlx_sram_chipsel_test.sv"
`include "nlx_sram_rstn_test.sv"

`endif//nlx_sram_TESTS_SVH

